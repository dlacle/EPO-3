configuration fa_behavioral_cfg of fa is
   for behavioral
   end for;
end fa_behavioral_cfg;
