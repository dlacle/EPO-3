configuration ha_behavioral_cfg of ha is
   for behavioral
   end for;
end ha_behavioral_cfg;
