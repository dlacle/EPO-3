library IEEE;
use IEEE.std_logic_1164.ALL;

entity shifter_right_tb is
end shifter_right_tb;



