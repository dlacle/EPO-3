configuration main_ytob_synthesised_cfg of main_ytob is
   for synthesised
   end for;
end main_ytob_synthesised_cfg;
