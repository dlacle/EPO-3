configuration zoomandposition_control_behavioural_cfg of zoomandposition_control is
   for behavioural
   end for;
end zoomandposition_control_behavioural_cfg;
