configuration main_seq_synthesised_cfg of main_seq is
   for synthesised
   end for;
end main_seq_synthesised_cfg;
