library IEEE;
use IEEE.std_logic_1164.ALL;

entity main_tb is
end main_tb;

