configuration shifter_left_2_behavioural_cfg of shifter_left_2 is
   for behavioural
   end for;
end shifter_left_2_behavioural_cfg;
