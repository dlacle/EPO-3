configuration ycounter_behavioural_cfg of ycounter is
   for behavioural
   end for;
end ycounter_behavioural_cfg;
