library IEEE;
use IEEE.std_logic_1164.ALL;

entity main_seq_tb is
end main_seq_tb;

