configuration register_a_structural_cfg of register_a is
   for structural
   end for;
end register_a_structural_cfg;
