library IEEE;
use IEEE.std_logic_1164.ALL;

entity shifter_right is
   port(s_in : in  std_logic_vector(11 downto 0);
	 s_out : out std_logic_vector(11 downto 0)
);
end shifter_right;

