configuration shifter_right_behavioural_cfg of shifter_right is
   for behavioural
   end for;
end shifter_right_behavioural_cfg;
