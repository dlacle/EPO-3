configuration unsignedto2_behaviour_cfg of unsignedto2 is
   for behaviour
   end for;
end unsignedto2_behaviour_cfg;
