configuration main_synthesised_cfg of main is
   for synthesised
   end for;
end main_synthesised_cfg;
