configuration main_xtoa_synthesised_cfg of main_xtoa is
   for synthesised
   end for;
end main_xtoa_synthesised_cfg;
