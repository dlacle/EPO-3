configuration main_ytobtb_behaviour_cfg of main_ytobtb is
   for behaviour
      for all: main_ytob use configuration work.main_ytob_synthesised_cfg;
      end for;
   end for;
end main_ytobtb_behaviour_cfg;
