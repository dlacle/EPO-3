configuration mux_position_behavioural_cfg of mux_position is
   for behavioural
   end for;
end mux_position_behavioural_cfg;
