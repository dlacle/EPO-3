configuration shifter_right_synthesised_cfg of shifter_right is
   for synthesised
   end for;
end shifter_right_synthesised_cfg;
